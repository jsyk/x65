/**
 * NORA Registers inside of the 0x9Fxx block.
 * This also instantiates all the requisite slaves. ????
 */
module regs
(
    // Global signals
    input           clk6x,      // 48MHz
    input           resetn,     // sync reset

);


endmodule